module OVERTURE (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_IOSwitch # (.UUID(64'd4 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_0 (.in(wire_1), .en(wire_22), .out(arch_output_value));
  TC_Splitter8 # (.UUID(64'd3075346555542787867 ^ UUID)) Splitter8_1 (.in(wire_4), .out0(wire_29), .out1(wire_33), .out2(wire_6), .out3(wire_11), .out4(wire_34), .out5(wire_19), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd2836361948119126518 ^ UUID)) Decoder3_2 (.dis(wire_26), .sel0(wire_29), .sel1(wire_33), .sel2(wire_6), .out0(wire_5), .out1(wire_8), .out2(wire_30), .out3(wire_25), .out4(wire_23), .out5(wire_20), .out6(wire_22), .out7());
  TC_Decoder3 # (.UUID(64'd1350450359641734825 ^ UUID)) Decoder3_3 (.dis(wire_26), .sel0(wire_11), .sel1(wire_34), .sel2(wire_19), .out0(wire_13), .out1(wire_0), .out2(wire_12), .out3(wire_28), .out4(wire_31), .out5(wire_32), .out6(wire_27), .out7());
  TC_Not # (.UUID(64'd2921486240680985383 ^ UUID), .BIT_WIDTH(64'd1)) Not_4 (.in(wire_10), .out(wire_26));
  TC_Switch # (.UUID(64'd4553160874405357450 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_5 (.en(wire_7), .in(wire_18), .out(wire_1_4));
  TC_Or # (.UUID(64'd2341608836636325000 ^ UUID), .BIT_WIDTH(64'd1)) Or_6 (.in0(wire_25), .in1(wire_7), .out(wire_16));
  TC_Switch # (.UUID(64'd888663386662975279 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_7 (.en(wire_27), .in(arch_input_value), .out(wire_1_5));
  TC_Counter # (.UUID(64'd2065154129327891408 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd1)) Counter8_8 (.clk(clk), .rst(rst), .save(wire_36), .in(wire_14), .out(wire_35));
  TC_Switch # (.UUID(64'd1906344177036918899 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_9 (.en(wire_9), .in(wire_4), .out(wire_1_0));
  TC_Or # (.UUID(64'd2414690846422019408 ^ UUID), .BIT_WIDTH(64'd1)) Or_10 (.in0(wire_5), .in1(wire_9), .out(wire_3));
  TC_Switch # (.UUID(64'd1109943128734162865 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_11 (.en(wire_17), .in(wire_15), .out(wire_36));
  TC_Program8_4 # (.UUID(64'd5 ^ UUID), .DEFAULT_FILE_NAME("Program8_4_5.w8.bin"), .ARG_SIG("Program8_4_5=%s")) Program8_4_12 (.clk(clk), .rst(rst), .address(wire_35), .out0(wire_4), .out1(), .out2(), .out3());
  DEC # (.UUID(64'd3584181306077434485 ^ UUID)) DEC_13 (.clk(clk), .rst(rst), .OPCODE(wire_4), .IMMEDIATE(wire_9), .CONDITION(wire_17), .CALCULATION(wire_7), .COPY(wire_10));
  ALUz_Compact # (.UUID(64'd3204575145873368728 ^ UUID)) ALUz_Compact_14 (.clk(clk), .rst(rst), .Code(wire_4), .Input_1(wire_24), .Input_2(wire_2), .Output(wire_18));
  CONDz_Compact # (.UUID(64'd1875835048430223602 ^ UUID)) CONDz_Compact_15 (.clk(clk), .rst(rst), .Condition(wire_4), .Input(wire_21), .Result(wire_15));
  RegisterPlus # (.UUID(64'd100000 ^ UUID)) RegisterPlus_16 (.clk(clk), .rst(rst), .Load(wire_13), .Save_value(wire_1), .Save(wire_3), .Always_output(wire_14), .Output(wire_1_1));
  RegisterPlus # (.UUID(64'd110000 ^ UUID)) RegisterPlus_17 (.clk(clk), .rst(rst), .Load(wire_0), .Save_value(wire_1), .Save(wire_8), .Always_output(wire_24), .Output(wire_1_2));
  RegisterPlus # (.UUID(64'd120000 ^ UUID)) RegisterPlus_18 (.clk(clk), .rst(rst), .Load(wire_12), .Save_value(wire_1), .Save(wire_30), .Always_output(wire_2), .Output(wire_1_3));
  RegisterPlus # (.UUID(64'd130000 ^ UUID)) RegisterPlus_19 (.clk(clk), .rst(rst), .Load(wire_28), .Save_value(wire_1), .Save(wire_16), .Always_output(wire_21), .Output(wire_1_6));
  RegisterPlus # (.UUID(64'd140000 ^ UUID)) RegisterPlus_20 (.clk(clk), .rst(rst), .Load(wire_31), .Save_value(wire_1), .Save(wire_23), .Always_output(), .Output(wire_1_7));
  RegisterPlus # (.UUID(64'd150000 ^ UUID)) RegisterPlus_21 (.clk(clk), .rst(rst), .Load(wire_32), .Save_value(wire_1), .Save(wire_20), .Always_output(), .Output(wire_1_8));

  wire [0:0] wire_0;
  wire [7:0] wire_1;
  wire [7:0] wire_1_0;
  wire [7:0] wire_1_1;
  wire [7:0] wire_1_2;
  wire [7:0] wire_1_3;
  wire [7:0] wire_1_4;
  wire [7:0] wire_1_5;
  wire [7:0] wire_1_6;
  wire [7:0] wire_1_7;
  wire [7:0] wire_1_8;
  assign wire_1 = wire_1_0|wire_1_1|wire_1_2|wire_1_3|wire_1_4|wire_1_5|wire_1_6|wire_1_7|wire_1_8;
  wire [7:0] wire_2;
  wire [0:0] wire_3;
  wire [7:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [7:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [7:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [7:0] wire_21;
  wire [0:0] wire_22;
  assign arch_output_enable = wire_22;
  wire [0:0] wire_23;
  wire [7:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  assign arch_input_enable = wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [7:0] wire_35;
  wire [0:0] wire_36;

endmodule
